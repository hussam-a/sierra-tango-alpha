module mux2_1(output2, x, y, sel);  wire _00_;  wire _01_;  wire _02_;  wire _03_;  wire _04_;  wire _05_;  wire _06_;  wire _07_;  output [3:0] output2;  input sel;  input [3:0] x;  input [3:0] y;  INVX1 _08_ (    .A(x[0]),    .Y(_00_)  );  NAND2X1 _09_ (    .A(y[0]),    .B(sel),    .Y(_01_)  );  OAI21X1 _10_ (    .A(sel),    .B(_00_),    .C(_01_),    .Y(output2[0])  );  INVX1 _11_ (    .A(x[1]),    .Y(_02_)  );  NAND2X1 _12_ (    .A(sel),    .B(y[1]),    .Y(_03_)  );  OAI21X1 _13_ (    .A(sel),    .B(_02_),    .C(_03_),    .Y(output2[1])  );  INVX1 _14_ (    .A(x[2]),    .Y(_04_)  );  NAND2X1 _15_ (    .A(sel),    .B(y[2]),    .Y(_05_)  );  OAI21X1 _16_ (    .A(sel),    .B(_04_),    .C(_05_),    .Y(output2[2])  );  INVX1 _17_ (    .A(x[3]),    .Y(_06_)  );  NAND2X1 _18_ (    .A(sel),    .B(y[3]),    .Y(_07_)  );  OAI21X1 _19_ (    .A(sel),    .B(_06_),    .C(_07_),    .Y(output2[3])  );endmodule
