module RtoR(clk, rst, a, b, f);  wire _0_;  wire _1_;  input a;  input b;  input clk;  wire comb2;  wire \dff1.D ;  wire \dff1.q ;  output f;  input rst;  INVX1 _2_ (    .A(a),    .Y(\dff1.D )  );  NAND2X1 _3_ (    .A(\dff1.q ),    .B(b),    .Y(comb2)  );  AND2X2 _4_ (    .A(\dff1.D ),    .B(rst),    .Y(_0_)  );  DFFPOSX1 _5_ (    .CLK(clk),    .D(_0_),    .Q(\dff1.q )  );  AND2X2 _6_ (    .A(comb2),    .B(rst),    .Y(_1_)  );  DFFPOSX1 _7_ (    .CLK(clk),    .D(_1_),    .Q(f)  );endmodule
