module mux4_1(output2, w, x, y, z, sel);  wire _00_;  wire _01_;  wire _02_;  wire _03_;  wire _04_;  wire _05_;  wire _06_;  wire _07_;  wire _08_;  wire _09_;  wire _10_;  wire _11_;  wire _12_;  wire _13_;  wire _14_;  wire _15_;  wire _16_;  wire _17_;  wire _18_;  wire _19_;  wire _20_;  wire _21_;  wire _22_;  wire _23_;  wire _24_;  wire _25_;  wire _26_;  wire _27_;  wire _28_;  wire _29_;  wire _30_;  wire _31_;  wire _32_;  wire _33_;  wire _34_;  wire _35_;  output [3:0] output2;  input [1:0] sel;  input [3:0] w;  input [3:0] x;  input [3:0] y;  input [3:0] z;  NAND2X1 _36_ (    .A(w[0]),    .B(_00_),    .Y(_01_)  );  INVX1 _37_ (    .A(sel[1]),    .Y(_02_)  );  INVX1 _38_ (    .A(z[0]),    .Y(_03_)  );  OAI21X1 _39_ (    .A(sel[0]),    .B(_02_),    .C(_03_),    .Y(_04_)  );  INVX1 _40_ (    .A(sel[0]),    .Y(_05_)  );  INVX1 _41_ (    .A(y[0]),    .Y(_06_)  );  NAND3X1 _42_ (    .A(sel[1]),    .B(_05_),    .C(_06_),    .Y(_07_)  );  AOI22X1 _43_ (    .A(_02_),    .B(sel[0]),    .C(_07_),    .D(_04_),    .Y(_08_)  );  AOI21X1 _44_ (    .A(sel[0]),    .B(x[0]),    .C(sel[1]),    .Y(_09_)  );  OAI21X1 _45_ (    .A(_09_),    .B(_08_),    .C(_01_),    .Y(output2[0])  );  NAND2X1 _46_ (    .A(w[1]),    .B(_00_),    .Y(_10_)  );  INVX1 _47_ (    .A(z[1]),    .Y(_11_)  );  NAND2X1 _48_ (    .A(sel[0]),    .B(_02_),    .Y(_12_)  );  NAND2X1 _49_ (    .A(sel[1]),    .B(_05_),    .Y(_13_)  );  NAND3X1 _50_ (    .A(_11_),    .B(_12_),    .C(_13_),    .Y(_14_)  );  INVX1 _51_ (    .A(y[1]),    .Y(_15_)  );  NAND3X1 _52_ (    .A(sel[1]),    .B(_05_),    .C(_15_),    .Y(_16_)  );  INVX1 _53_ (    .A(x[1]),    .Y(_17_)  );  OAI21X1 _54_ (    .A(_05_),    .B(_17_),    .C(_02_),    .Y(_18_)  );  NAND3X1 _55_ (    .A(_16_),    .B(_18_),    .C(_14_),    .Y(_19_)  );  NAND2X1 _56_ (    .A(_10_),    .B(_19_),    .Y(output2[1])  );  NAND2X1 _57_ (    .A(w[2]),    .B(_00_),    .Y(_20_)  );  INVX1 _58_ (    .A(z[2]),    .Y(_21_)  );  NAND3X1 _59_ (    .A(_21_),    .B(_12_),    .C(_13_),    .Y(_22_)  );  INVX1 _60_ (    .A(y[2]),    .Y(_23_)  );  NAND3X1 _61_ (    .A(sel[1]),    .B(_05_),    .C(_23_),    .Y(_24_)  );  INVX1 _62_ (    .A(x[2]),    .Y(_25_)  );  OAI21X1 _63_ (    .A(_05_),    .B(_25_),    .C(_02_),    .Y(_26_)  );  NAND3X1 _64_ (    .A(_24_),    .B(_26_),    .C(_22_),    .Y(_27_)  );  NAND2X1 _65_ (    .A(_20_),    .B(_27_),    .Y(output2[2])  );  NAND2X1 _66_ (    .A(w[3]),    .B(_00_),    .Y(_28_)  );  INVX1 _67_ (    .A(z[3]),    .Y(_29_)  );  NAND3X1 _68_ (    .A(_29_),    .B(_12_),    .C(_13_),    .Y(_30_)  );  INVX1 _69_ (    .A(y[3]),    .Y(_31_)  );  NAND3X1 _70_ (    .A(sel[1]),    .B(_05_),    .C(_31_),    .Y(_32_)  );  INVX1 _71_ (    .A(x[3]),    .Y(_33_)  );  OAI21X1 _72_ (    .A(_05_),    .B(_33_),    .C(_02_),    .Y(_34_)  );  NAND3X1 _73_ (    .A(_32_),    .B(_34_),    .C(_30_),    .Y(_35_)  );  NAND2X1 _74_ (    .A(_28_),    .B(_35_),    .Y(output2[3])  );  NOR2X1 _75_ (    .A(sel[1]),    .B(sel[0]),    .Y(_00_)  );endmodule
