module simpleR_R(a, d, clk, rst, y);  wire _0_;  wire _1_;  input a;  wire c;  input clk;  input d;  wire \dff2.D ;  input rst;  output y;  OR2X2 _2_ (    .A(c),    .B(a),    .Y(\dff2.D )  );  AND2X2 _3_ (    .A(d),    .B(rst),    .Y(_0_)  );  DFFPOSX1 _4_ (    .CLK(clk),    .D(_0_),    .Q(c)  );  AND2X2 _5_ (    .A(\dff2.D ),    .B(rst),    .Y(_1_)  );  DFFPOSX1 _6_ (    .CLK(clk),    .D(_1_),    .Q(y)  );endmodule
