module fourbitmux2X1ToRegToReg(out, x, y, sel, clk);  wire _00_;  wire _01_;  wire _02_;  wire _03_;  wire _04_;  wire _05_;  wire _06_;  wire _07_;  wire [3:0] \_mux4_1.out ;  input clk;  output [3:0] out;  wire [3:0] r1;  input sel;  input [3:0] x;  input [3:0] y;  DFFPOSX1 _08_ (    .CLK(clk),    .D(r1[0]),    .Q(out[0])  );  DFFPOSX1 _09_ (    .CLK(clk),    .D(r1[1]),    .Q(out[1])  );  DFFPOSX1 _10_ (    .CLK(clk),    .D(r1[2]),    .Q(out[2])  );  DFFPOSX1 _11_ (    .CLK(clk),    .D(r1[3]),    .Q(out[3])  );  DFFPOSX1 _12_ (    .CLK(clk),    .D(\_mux4_1.out [0]),    .Q(r1[0])  );  DFFPOSX1 _13_ (    .CLK(clk),    .D(\_mux4_1.out [1]),    .Q(r1[1])  );  DFFPOSX1 _14_ (    .CLK(clk),    .D(\_mux4_1.out [2]),    .Q(r1[2])  );  DFFPOSX1 _15_ (    .CLK(clk),    .D(\_mux4_1.out [3]),    .Q(r1[3])  );  INVX1 _16_ (    .A(x[0]),    .Y(_00_)  );  NAND2X1 _17_ (    .A(y[0]),    .B(sel),    .Y(_01_)  );  OAI21X1 _18_ (    .A(sel),    .B(_00_),    .C(_01_),    .Y(\_mux4_1.out [0])  );  INVX1 _19_ (    .A(x[1]),    .Y(_02_)  );  NAND2X1 _20_ (    .A(sel),    .B(y[1]),    .Y(_03_)  );  OAI21X1 _21_ (    .A(sel),    .B(_02_),    .C(_03_),    .Y(\_mux4_1.out [1])  );  INVX1 _22_ (    .A(x[2]),    .Y(_04_)  );  NAND2X1 _23_ (    .A(sel),    .B(y[2]),    .Y(_05_)  );  OAI21X1 _24_ (    .A(sel),    .B(_04_),    .C(_05_),    .Y(\_mux4_1.out [2])  );  INVX1 _25_ (    .A(x[3]),    .Y(_06_)  );  NAND2X1 _26_ (    .A(sel),    .B(y[3]),    .Y(_07_)  );  OAI21X1 _27_ (    .A(sel),    .B(_06_),    .C(_07_),    .Y(\_mux4_1.out [3])  );endmodule
